module bin2gray (
    
);
    
endmodule